module datapath(
    input wire clock, clear, 
    

)