module ripplecarryadder(
    input [31:0] A,B,
    output reg [31:0] CC,
    input wire Select
);
